----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    20:38:15 11/27/2016 
-- Design Name: 
-- Module Name:    mux2x1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux2x1 is
    Port ( A : in  STD_LOGIC_vector(7 downto 0);
           B : in  STD_LOGIC_vector(7 downto 0);
           sel : in  STD_LOGIC;
           output : out  STD_LOGIC_vector(7 downto 0));
end mux2x1;

architecture Behavioral of mux2x1 is

begin

with sel select output <=
   A when '0',
	B when '1',
	"XXXXXXXX" when others;


end Behavioral;

